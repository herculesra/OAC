CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
290 50 10 200 9
48 106 1872 1004
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
54 C:\Users\H�rcules\Desktop\Circuito Maker\CM60S\BOM.DAT
0 7
48 106 1872 1004
210763794 0
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 606 253 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
5 CLOCK
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 608 207 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 -16 9 -8
5 INPUT
-16 -26 19 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 721 170 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 801 170 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 895 167 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 977 167 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 Q0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
12 D Flip-Flop~
219 679 244 0 4 9
0 6 5 8 4
0
0 0 4208 0
3 DFF
-10 -53 11 -45
2 A1
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9914 0 0
0
0
12 D Flip-Flop~
219 763 244 0 4 9
0 4 5 9 3
0
0 0 4208 0
3 DFF
-10 -53 11 -45
2 A2
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3747 0 0
0
0
12 D Flip-Flop~
219 848 244 0 4 9
0 3 5 10 2
0
0 0 4208 0
3 DFF
-10 -53 11 -45
2 A3
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3549 0 0
0
0
12 D Flip-Flop~
219 947 244 0 4 9
0 2 5 11 7
0
0 0 4208 0
3 DFF
-10 -53 11 -45
2 A4
-7 -63 7 -55
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
7931 0 0
0
0
12
0 1 2 0 0 4096 0 0 5 2 0 2
895 208
895 185
4 1 2 0 0 4224 0 9 10 0 0 2
872 208
923 208
0 1 3 0 0 8192 0 0 4 4 0 3
803 208
801 208
801 188
4 1 3 0 0 4224 0 8 9 0 0 2
787 208
824 208
0 1 4 0 0 8192 0 0 3 6 0 3
720 208
721 208
721 188
4 1 4 0 0 4224 0 7 8 0 0 2
703 208
739 208
2 0 5 0 0 4096 0 7 0 0 10 2
655 226
655 253
2 0 5 0 0 0 0 8 0 0 10 2
739 226
739 253
2 0 5 0 0 0 0 9 0 0 10 2
824 226
824 253
1 2 5 0 0 4224 0 1 10 0 0 3
618 253
923 253
923 226
1 1 6 0 0 8320 0 2 7 0 0 3
620 207
620 208
655 208
4 1 7 0 0 8320 0 10 6 0 0 3
971 208
977 208
977 185
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
