CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 9
0 71 1920 1040
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
54 C:\Users\H�rcules\Desktop\Circuito Maker\CM60S\BOM.DAT
0 7
0 71 1920 1040
143655186 0
0
6 Title:
5 Name:
0
0
0
8
13 Logic Switch~
5 528 167 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-10 15 4 23
1 A
-5 -23 2 -15
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 537 301 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-5 18 9 26
1 B
-2 -30 5 -22
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
14 Logic Display~
6 863 275 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 857 157 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6153 0 0
0
0
9 Inverter~
13 616 302 0 2 22
0 3 8
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 2 3 0
1 U
5394 0 0
0
0
9 Inverter~
13 592 164 0 2 22
0 4 7
0
0 0 112 0
6 74LS04
-21 -19 21 -11
0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
15

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0
65 0 0 0 6 1 3 0
1 U
7734 0 0
0
0
10 2-In NAND~
219 735 293 0 3 22
0 6 8 5
0
0 0 112 0
4 7400
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
10 2-In NAND~
219 730 175 0 3 22
0 7 5 6
0
0 0 112 0
4 7400
-7 -24 21 -16
0
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 -1766218101
65 0 0 0 4 1 2 0
1 U
3747 0 0
0
0
8
1 1 3 0 0 8320 0 2 5 0 0 3
549 301
549 302
601 302
1 1 4 0 0 4224 0 1 6 0 0 4
540 167
555 167
555 164
577 164
1 0 5 0 0 4224 0 3 0 0 8 2
863 293
815 293
1 0 6 0 0 8320 0 4 0 0 7 3
857 175
857 177
845 177
2 1 7 0 0 12416 0 6 8 0 0 4
613 164
650 164
650 166
706 166
2 2 8 0 0 4224 0 5 7 0 0 2
637 302
711 302
3 1 6 0 0 16512 0 8 7 0 0 7
757 175
757 177
845 177
845 212
683 212
683 284
711 284
3 2 5 0 0 12416 0 7 8 0 0 6
762 293
815 293
815 250
694 250
694 184
706 184
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-006 1e-007 1e-007
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
